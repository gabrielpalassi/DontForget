LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY mux_8x1_n IS
    GENERIC (
        CONSTANT BITS : INTEGER := 4
    );
    PORT (
        D0 : IN STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0);
        D1 : IN STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0);
        D2 : IN STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0);
        D3 : IN STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0);
        D4 : IN STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0);
        D5 : IN STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0);
        D6 : IN STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0);
        D7 : IN STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0);
        SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
        MUX_OUT : OUT STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE behav OF mux_8x1_n IS
BEGIN
    MUX_OUT <= D7 WHEN (SEL = "111") ELSE
        D6 WHEN (SEL = "110") ELSE
        D5 WHEN (SEL = "101") ELSE
        D4 WHEN (SEL = "100") ELSE
        D3 WHEN (SEL = "011") ELSE
        D2 WHEN (SEL = "010") ELSE
        D1 WHEN (SEL = "001") ELSE
        D0 WHEN (SEL = "000") ELSE
        (OTHERS => '1');
END ARCHITECTURE behav;